library verilog;
use verilog.vl_types.all;
entity ise_proj_vlg_vec_tst is
end ise_proj_vlg_vec_tst;
