
//------> ./rtl_mgc_ioport.v 
//------------------------------------------------------------------
//                M G C _ I O P O R T _ C O M P S
//------------------------------------------------------------------

//------------------------------------------------------------------
//                       M O D U L E S
//------------------------------------------------------------------

//------------------------------------------------------------------
//-- INPUT ENTITIES
//------------------------------------------------------------------

module mgc_in_wire (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output [width-1:0] d;
  output             lz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule
//------------------------------------------------------------------

module mgc_chan_in (ld, vd, d, lz, vz, z, size, req_size, sizez, sizelz);

  parameter integer rscid = 1;
  parameter integer width = 8;
  parameter integer sz_width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;
  output [sz_width-1:0] size;
  input              req_size;
  input  [sz_width-1:0] sizez;
  output             sizelz;


  wire               vd;
  wire   [width-1:0] d;
  wire               lz;
  wire   [sz_width-1:0] size;
  wire               sizelz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;
  assign size = sizez;
  assign sizelz = req_size;

endmodule


//------------------------------------------------------------------
//-- OUTPUT ENTITIES
//------------------------------------------------------------------

module mgc_out_stdreg (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  input  [width-1:0] d;
  output             lz;
  output [width-1:0] z;

  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_out_prereg_en (ld, d, lz, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    wire               lz;
    wire   [width-1:0] z;

    assign z = d;
    assign lz = ld;

endmodule

//------------------------------------------------------------------
//-- INOUT ENTITIES
//------------------------------------------------------------------

module mgc_inout_stdreg_en (ldin, din, ldout, dout, lzin, lzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    output             lzin;
    output             lzout;
    inout  [width-1:0] z;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign z = ldout ? dout : {width{1'bz}};

endmodule

//------------------------------------------------------------------
module hid_tribuf( I_SIG, ENABLE, O_SIG);
  parameter integer width = 8;

  input [width-1:0] I_SIG;
  input ENABLE;
  inout [width-1:0] O_SIG;

  assign O_SIG = (ENABLE) ? I_SIG : { width{1'bz}};

endmodule
//------------------------------------------------------------------

module mgc_inout_stdreg_wait (ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;
    wire   ldout_and_vzout;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign vdout = vzout ;
    assign ldout_and_vzout = ldout && vzout ;

    hid_tribuf #(width) tb( .I_SIG(dout),
                            .ENABLE(ldout_and_vzout),
                            .O_SIG(z) );

endmodule

//------------------------------------------------------------------

module mgc_inout_buf_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    hid_tribuf #(width) tb( .I_SIG(z_buf),
                            .ENABLE((lzout_buf && (!ldin) && vzout) ),
                            .O_SIG(z)  );

    mgc_out_buf_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFF
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );


endmodule

module mgc_inout_fifo_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer ph_log2 = 3;     // log2(fifo_sz)
    parameter integer pwropt  = 0;     // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               comb;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    assign comb = (lzout_buf && (!ldin) && vzout);

    hid_tribuf #(width) tb2( .I_SIG(z_buf), .ENABLE(comb), .O_SIG(z)  );

    mgc_out_fifo_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
    )
    FIFO
    (
        .clk   (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );

endmodule

//------------------------------------------------------------------
//-- I/O SYNCHRONIZATION ENTITIES
//------------------------------------------------------------------

module mgc_io_sync (ld, lz);

    input  ld;
    output lz;

    assign lz = ld;

endmodule

module mgc_bsync_rdy (rd, rz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 0;

    input  rd;
    output rz;

    wire   rz;

    assign rz = rd;

endmodule

module mgc_bsync_vld (vd, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 0;
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule

module mgc_bsync_rv (rd, vd, rz, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 1;

    input  rd;
    output vd;
    output rz;
    input  vz;

    wire   vd;
    wire   rz;

    assign rz = rd;
    assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_sync (ldin, vdin, ldout, vdout);

  input  ldin;
  output vdin;
  input  ldout;
  output vdout;

  wire   vdin;
  wire   vdout;

  assign vdin = ldout;
  assign vdout = ldin;

endmodule

///////////////////////////////////////////////////////////////////////////////
// dummy function used to preserve funccalls for modulario
// it looks like a memory read to the caller
///////////////////////////////////////////////////////////////////////////////
module funccall_inout (d, ad, bd, z, az, bz);

  parameter integer ram_id = 1;
  parameter integer width = 8;
  parameter integer addr_width = 8;

  output [width-1:0]       d;
  input  [addr_width-1:0]  ad;
  input                    bd;
  input  [width-1:0]       z;
  output [addr_width-1:0]  az;
  output                   bz;

  wire   [width-1:0]       d;
  wire   [addr_width-1:0]  az;
  wire                     bz;

  assign d  = z;
  assign az = ad;
  assign bz = bd;

endmodule


///////////////////////////////////////////////////////////////////////////////
// inlinable modular io not otherwise found in mgc_ioport
///////////////////////////////////////////////////////////////////////////////

module modulario_en_in (vd, d, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output             vd;
  output [width-1:0] d;
  input              vz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               vd;

  assign d = z;
  assign vd = vz;

endmodule

//------> ./rtl_mgc_ioport_v2001.v 
//------------------------------------------------------------------

module mgc_out_reg_pos (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(posedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(posedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg_neg (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(negedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(negedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg (clk, en, arst, srst, ld, d, lz, z); // Not Supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;


    generate
    if (ph_clk == 1'b0)
    begin: NEG_EDGE

        mgc_out_reg_neg
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_neg_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    else
    begin: POS_EDGE

        mgc_out_reg_pos
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_pos_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    endgenerate

endmodule




//------------------------------------------------------------------

module mgc_out_buf_wait (clk, en, arst, srst, ld, vd, d, vz, lz, z); // Not supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    output             vd;
    input  [width-1:0] d;
    output             lz;
    input              vz;
    output [width-1:0] z;

    wire               filled;
    wire               filled_next;
    wire   [width-1:0] abuf;
    wire               lbuf;


    assign filled_next = (filled & (~vz)) | (filled & ld) | (ld & (~vz));

    assign lbuf = ld & ~(filled ^ vz);

    assign vd = vz | ~filled;

    assign lz = ld | filled;

    assign z = (filled) ? abuf : d;

    wire dummy;
    wire dummy_bufreg_lz;

    // Output registers:
    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (1'b1),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    STATREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (filled_next),
        .d       (1'b0),       // input d is unused
        .lz      (filled),
        .z       (dummy)            // output z is unused
    );

    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (lbuf),
        .d       (d),
        .lz      (dummy_bufreg_lz),
        .z       (abuf)
    );

endmodule

//------------------------------------------------------------------

module mgc_out_fifo_wait (clk, en, arst, srst, ld, vd, d, lz, vz,  z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1; // clock enable polarity
    parameter         ph_arst = 1'b1; // async reset polarity
    parameter         ph_srst = 1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt


    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;

    wire    [31:0]      size;


      // Output registers:
 mgc_out_fifo_wait_core#(
        .rscid   (rscid),
        .width   (width),
        .sz_width (32),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
        ) CORE (
        .clk (clk),
        .en (en),
        .arst (arst),
        .srst (srst),
        .ld (ld),
        .vd (vd),
        .d (d),
        .lz (lz),
        .vz (vz),
        .z (z),
        .size (size)
        );

endmodule



module mgc_out_fifo_wait_core (clk, en, arst, srst, ld, vd, d, lz, vz,  z, size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt

   localparam integer  fifo_b = width * fifo_sz;

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;
    output    [sz_width-1:0]      size;

    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat_pre;
    wire     [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] en_l;
    reg      [(((fifo_sz > 0) ? fifo_sz : 1)-1)/8:0] en_l_s;

    reg       [width-1:0] buff_nxt;

    reg                   stat_nxt;
    reg                   stat_before;
    reg                   stat_after;
    reg                   en_l_var;

    integer               i;
    genvar                eni;

    wire [32:0]           size_t;
    reg [31:0]            count;
    reg [31:0]            count_t;
    reg [32:0]            n_elem;
// pragma translate_off
    reg [31:0]            peak;
// pragma translate_on

    wire [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] dummy_statreg_lz;
    wire [( (fifo_b > 0) ? fifo_b : 1)-1:0] dummy_bufreg_lz;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = (count - (vz && stat[fifo_sz-1])) + ld;
      assign size = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          if (i != 0)
            stat_before = stat[i-1];
          else
            stat_before = 1'b0;

          if (i != (fifo_sz-1))
            stat_after = stat[i+1];
          else
            stat_after = 1'b1;

          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));

          stat_pre[i] = stat_nxt;
          en_l_var = 1'b1;
          if (!stat_nxt)
            begin
              buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end
          else if (vz && stat_before)
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
          else if (ld && !((vz && stat_before) || ((!vz) && stat[i])))
            buff_nxt = d;
          else
            begin
              if (pwropt == 0)
                buff_nxt[0+:width] = buff[width*i+:width];
              else
                buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if ((stat_after == 1'b1) && (stat[i] == 1'b0))
            n_elem = ($unsigned(fifo_sz) - 1) - i;
        end

        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b1;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b0;

        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if ((i%'d2) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]|stat_pre[i-1]);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]|stat_pre[i-1]);
          end
        end

        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = { {(32-ph_log2){1'b0}}, fifo_sz};
        else
          count_t = n_elem[31:0];
        count = count_t;
// pragma translate_off
        if ( peak < count )
          peak = count;
// pragma translate_on
      end

      if (pwropt == 0)
      begin: NOCGFIFO
        // Output registers:
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        STATREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
        );
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_b),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        BUFREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre),
            .lz      (dummy_bufreg_lz[0]),
            .z       (buff)
        );
      end
      else
      begin: CGFIFO
        // Output registers:
        if ( pwropt > 1)
        begin: CGSTATFIFO2
          for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
          begin: pwroptGEN1
            mgc_out_reg
            #(
              .rscid   (rscid),
              .width   (1),
              .ph_clk  (ph_clk),
              .ph_en   (ph_en),
              .ph_arst (ph_arst),
              .ph_srst (ph_srst)
            )
            STATREG
            (
              .clk     (clk),
              .en      (en_l_s[eni/8]),
              .arst    (arst),
              .srst    (srst),
              .ld      (1'b1),
              .d       (stat_pre[eni]),
              .lz      (dummy_statreg_lz[eni]),
              .z       (stat[eni])
            );
          end
        end
        else
        begin: CGSTATFIFO
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          STATREG
          (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
          );
        end
        for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
        begin: pwroptGEN2
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (width),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          BUFREG
          (
            .clk     (clk),
            .en      (en_l[eni]),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre[width*eni+:width]),
            .lz      (dummy_bufreg_lz[eni]),
            .z       (buff[width*eni+:width])
          );
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign size = ld && !vz;
    end
    endgenerate

endmodule

//------------------------------------------------------------------
//-- PIPE ENTITIES
//------------------------------------------------------------------
/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 */
// two clock pipe
module mgc_pipe (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, size, req_size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer pwropt  = 0; // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output [sz_width-1:0]      size;
    input              req_size;


    mgc_out_fifo_wait_core
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz),
        .pwropt   (pwropt)
    )
    FIFO
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (vdin),
        .vz      (ldin),
        .z       (din),
        .size    (size)
    );

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2011a.126 Production Release
//  HLS Date:       Wed Aug  8 00:52:07 PDT 2012
// 
//  Generated by:   oh1015@EEWS104A-006
//  Generated date: Tue Mar 08 14:56:50 2016
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    mean_vga_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module mean_vga_core_fsm (
  clk, rst, fsm_output, st_SHIFT_tr0, st_FRAME_2_tr0
);
  input clk;
  input rst;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;
  input st_SHIFT_tr0;
  input st_FRAME_2_tr0;


  // FSM State Type Declaration for mean_vga_core_fsm_1
  parameter
    st_main = 3'd0,
    st_FRAME = 3'd1,
    st_SHIFT = 3'd2,
    st_FRAME_1 = 3'd3,
    st_FRAME_2 = 3'd4,
    state_x = 3'b000;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : mean_vga_core_fsm_1
    case (state_var)
      st_main : begin
        fsm_output = 5'b1;
        state_var_NS = st_FRAME;
      end
      st_FRAME : begin
        fsm_output = 5'b10;
        state_var_NS = st_SHIFT;
      end
      st_SHIFT : begin
        fsm_output = 5'b100;
        if ( st_SHIFT_tr0 ) begin
          state_var_NS = st_FRAME_1;
        end
        else begin
          state_var_NS = st_SHIFT;
        end
      end
      st_FRAME_1 : begin
        fsm_output = 5'b1000;
        state_var_NS = st_FRAME_2;
      end
      st_FRAME_2 : begin
        fsm_output = 5'b10000;
        if ( st_FRAME_2_tr0 ) begin
          state_var_NS = st_main;
        end
        else begin
          state_var_NS = st_FRAME;
        end
      end
      default : begin
        fsm_output = 5'b00000;
        state_var_NS = st_main;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= st_main;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mean_vga_core
// ------------------------------------------------------------------


module mean_vga_core (
  clk, rst, vin_rsc_mgc_in_wire_d, vout_rsc_mgc_out_stdreg_d
);
  input clk;
  input rst;
  input [749:0] vin_rsc_mgc_in_wire_d;
  output [149:0] vout_rsc_mgc_out_stdreg_d;
  reg [149:0] vout_rsc_mgc_out_stdreg_d;


  // Interconnect Declarations
  wire [4:0] fsm_output;
  reg [29:0] regs_regs_0_1_lpi_2;
  reg [5:0] io_read_vout_rsc_d_sdt_sg1_lpi_2;
  reg [3:0] io_read_vout_rsc_d_sdt_sg2_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_1_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg3_lpi_2;
  reg [5:0] io_read_vout_rsc_d_sdt_sg5_lpi_2;
  reg [3:0] io_read_vout_rsc_d_sdt_sg6_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg4_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg7_lpi_2;
  reg [5:0] io_read_vout_rsc_d_sdt_sg9_lpi_2;
  reg [3:0] io_read_vout_rsc_d_sdt_sg10_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg8_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg11_lpi_2;
  reg [5:0] io_read_vout_rsc_d_sdt_sg13_lpi_2;
  reg [3:0] io_read_vout_rsc_d_sdt_sg14_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg12_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg15_lpi_2;
  reg [5:0] io_read_vout_rsc_d_sdt_sg17_lpi_2;
  reg [3:0] io_read_vout_rsc_d_sdt_sg18_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg16_lpi_2;
  reg [9:0] io_read_vout_rsc_d_sdt_sg19_lpi_2;
  reg [2:0] FRAME_p_1_sva;
  reg [29:0] regs_regs_0_1_lpi_3;
  reg [29:0] regs_operator_din_1_sva;
  reg [29:0] regs_regs_0_1_lpi_3_dfm;
  reg equal_tmp;
  reg equal_tmp_1;
  reg equal_tmp_2;
  reg equal_tmp_3;
  reg [9:0] io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm;
  reg [3:0] io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm;
  reg [5:0] io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm;
  reg [3:0] io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm;
  reg [5:0] io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm;
  reg [3:0] io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm;
  reg [5:0] io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm;
  reg [3:0] io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm;
  reg [5:0] io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm;
  reg [3:0] io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm;
  reg [5:0] io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm;
  reg [9:0] io_read_vout_rsc_d_sdt_1_lpi_2_dfm;
  reg [2:0] FRAME_p_1_sva_1;
  reg FRAME_slc_itm;
  reg SHIFT_i_1_sva_2_sg1;
  reg [1:0] SHIFT_i_1_sva_3;
  wire and_13_cse;
  wire nor_9_cse;
  wire nor_7_cse;
  wire nor_8_cse;
  wire [11:0] FRAME_acc_7_psp_sva;
  wire [12:0] nl_FRAME_acc_7_psp_sva;
  wire [3:0] z_out;
  wire [4:0] nl_z_out;
  wire [9:0] io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm_mx0;
  wire [3:0] io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm_mx0;
  wire [5:0] io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm_mx0;
  wire [3:0] io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm_mx0;
  wire [5:0] io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm_mx0;
  wire [3:0] io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm_mx0;
  wire [5:0] io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm_mx0;
  wire [3:0] io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm_mx0;
  wire [5:0] io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm_mx0;
  wire [3:0] io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm_mx0;
  wire [5:0] io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm_mx0;
  wire [9:0] io_read_vout_rsc_d_sdt_1_lpi_2_dfm_mx0;
  wire [5:0] FRAME_or_3_psp_sva;
  wire [9:0] FRAME_or_psp_sva;
  wire [11:0] FRAME_acc_6_psp_sva;
  wire [12:0] nl_FRAME_acc_6_psp_sva;
  wire [2:0] acc_imod_1_sva;
  wire [3:0] nl_acc_imod_1_sva;
  wire [3:0] acc_1_psp_sva;
  wire [4:0] nl_acc_1_psp_sva;
  wire or_161_tmp;
  wire and_cse;
  wire and_34_cse;

  wire[2:0] mux_47_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_mean_vga_core_fsm_inst_st_SHIFT_tr0;
  assign nl_mean_vga_core_fsm_inst_st_SHIFT_tr0 = z_out[2];
  wire [0:0] nl_mean_vga_core_fsm_inst_st_FRAME_2_tr0;
  assign nl_mean_vga_core_fsm_inst_st_FRAME_2_tr0 = ~ FRAME_slc_itm;
  mean_vga_core_fsm mean_vga_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .st_SHIFT_tr0(nl_mean_vga_core_fsm_inst_st_SHIFT_tr0),
      .st_FRAME_2_tr0(nl_mean_vga_core_fsm_inst_st_FRAME_2_tr0)
    );
  assign or_161_tmp = (SHIFT_i_1_sva_3[0]) | (SHIFT_i_1_sva_3[1]) | SHIFT_i_1_sva_2_sg1;
  assign and_cse = (~ or_161_tmp) & (fsm_output[2]);
  assign and_34_cse = or_161_tmp & (fsm_output[2]);
  assign nor_9_cse = ~((FRAME_p_1_sva[1]) | (FRAME_p_1_sva[0]));
  assign nor_7_cse = ~((FRAME_p_1_sva[2]) | (FRAME_p_1_sva[1]));
  assign nor_8_cse = ~((FRAME_p_1_sva[2]) | (FRAME_p_1_sva[0]));
  assign io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg19_lpi_2
      , FRAME_or_psp_sva}, equal_tmp_3);
  assign io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm_mx0 = MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg18_lpi_2
      , (FRAME_acc_7_psp_sva[9:6])}, equal_tmp_3);
  assign io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm_mx0 = MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg17_lpi_2
      , FRAME_or_3_psp_sva}, equal_tmp_3);
  assign io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg16_lpi_2
      , (FRAME_acc_7_psp_sva[9:0])}, equal_tmp_3);
  assign io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg15_lpi_2
      , FRAME_or_psp_sva}, equal_tmp_2);
  assign io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm_mx0 = MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg14_lpi_2
      , (FRAME_acc_7_psp_sva[9:6])}, equal_tmp_2);
  assign io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm_mx0 = MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg13_lpi_2
      , FRAME_or_3_psp_sva}, equal_tmp_2);
  assign io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg12_lpi_2
      , (FRAME_acc_7_psp_sva[9:0])}, equal_tmp_2);
  assign io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg11_lpi_2
      , FRAME_or_psp_sva}, equal_tmp_1);
  assign io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm_mx0 = MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg10_lpi_2
      , (FRAME_acc_7_psp_sva[9:6])}, equal_tmp_1);
  assign io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm_mx0 = MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg9_lpi_2
      , FRAME_or_3_psp_sva}, equal_tmp_1);
  assign io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg8_lpi_2
      , (FRAME_acc_7_psp_sva[9:0])}, equal_tmp_1);
  assign io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg7_lpi_2
      , FRAME_or_psp_sva}, equal_tmp);
  assign io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm_mx0 = MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg6_lpi_2
      , (FRAME_acc_7_psp_sva[9:6])}, equal_tmp);
  assign io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm_mx0 = MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg5_lpi_2
      , FRAME_or_3_psp_sva}, equal_tmp);
  assign io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg4_lpi_2
      , (FRAME_acc_7_psp_sva[9:0])}, equal_tmp);
  assign io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg3_lpi_2
      , FRAME_or_psp_sva}, and_13_cse);
  assign io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm_mx0 = MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg2_lpi_2
      , (FRAME_acc_7_psp_sva[9:6])}, and_13_cse);
  assign io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm_mx0 = MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg1_lpi_2
      , FRAME_or_3_psp_sva}, and_13_cse);
  assign io_read_vout_rsc_d_sdt_1_lpi_2_dfm_mx0 = MUX_v_10_2_2({io_read_vout_rsc_d_sdt_1_lpi_2
      , (FRAME_acc_7_psp_sva[9:0])}, and_13_cse);
  assign nl_FRAME_acc_7_psp_sva = conv_u2s_10_12({(FRAME_acc_6_psp_sva[11]) , (conv_u2u_8_9({(FRAME_acc_6_psp_sva[11])
      , 1'b0 , (FRAME_acc_6_psp_sva[11]) , 1'b0 , (FRAME_acc_6_psp_sva[11]) , 1'b0
      , (signext_2_1(FRAME_acc_6_psp_sva[7]))}) + conv_u2u_8_9(readslicef_9_8_1((({(FRAME_acc_6_psp_sva[9])
      , 1'b0 , (FRAME_acc_6_psp_sva[9]) , 1'b0 , (FRAME_acc_6_psp_sva[9]) , 1'b0
      , (signext_2_1(FRAME_acc_6_psp_sva[5])) , 1'b1}) + conv_u2u_8_9({(readslicef_8_7_1((conv_u2u_7_8({(FRAME_acc_6_psp_sva[7])
      , 1'b0 , (FRAME_acc_6_psp_sva[5]) , 1'b0 , (signext_2_1(FRAME_acc_6_psp_sva[9]))
      , 1'b1}) + conv_u2u_6_8({(FRAME_acc_6_psp_sva[6]) , 1'b0 , (FRAME_acc_6_psp_sva[6])
      , 1'b0 , (FRAME_acc_6_psp_sva[6]) , (acc_imod_1_sva[1])})))) , (~ (readslicef_3_1_2((({1'b1
      , (acc_imod_1_sva[0]) , 1'b1}) + conv_u2s_2_3({(~ (acc_imod_1_sva[1])) , (~
      (acc_imod_1_sva[2]))})))))})))))}) + conv_s2s_10_12(conv_u2s_9_10({(FRAME_acc_6_psp_sva[10])
      , 1'b0 , (FRAME_acc_6_psp_sva[10]) , 1'b0 , (FRAME_acc_6_psp_sva[10]) , 1'b0
      , (FRAME_acc_6_psp_sva[10]) , 1'b0 , (FRAME_acc_6_psp_sva[10])}) + conv_s2s_8_10(readslicef_9_8_1((conv_u2s_8_9({(FRAME_acc_6_psp_sva[8])
      , 1'b0 , (FRAME_acc_6_psp_sva[8]) , 1'b0 , (FRAME_acc_6_psp_sva[8]) , 1'b0
      , (FRAME_acc_6_psp_sva[8]) , 1'b1}) + conv_s2s_7_9({(readslicef_7_6_1((conv_s2s_5_7({(readslicef_5_4_1((conv_s2s_4_5({(readslicef_4_3_1((conv_u2s_3_4({(FRAME_acc_6_psp_sva[3])
      , (FRAME_acc_6_psp_sva[1]) , 1'b1}) + conv_s2s_3_4({1'b1 , (FRAME_acc_6_psp_sva[2])
      , (FRAME_acc_6_psp_sva[3])})))) , 1'b1}) + conv_s2s_3_5({(acc_1_psp_sva[3:2])
      , (FRAME_acc_6_psp_sva[4])})))) , 1'b1}) + conv_u2s_5_7({(FRAME_acc_6_psp_sva[7])
      , (FRAME_acc_6_psp_sva[4]) , (signext_2_1(FRAME_acc_6_psp_sva[11])) , (acc_1_psp_sva[1])}))))
      , (~ (acc_imod_1_sva[2]))})))));
  assign FRAME_acc_7_psp_sva = nl_FRAME_acc_7_psp_sva[11:0];
  assign FRAME_or_3_psp_sva = (FRAME_acc_7_psp_sva[5:0]) | (signext_6_2(FRAME_acc_7_psp_sva[11:10]));
  assign FRAME_or_psp_sva = (FRAME_acc_7_psp_sva[9:0]) | ({4'b0 , (signext_6_2(FRAME_acc_7_psp_sva[11:10]))});
  assign nl_FRAME_acc_6_psp_sva = conv_u2u_11_12(conv_u2u_10_11(regs_regs_0_1_lpi_3_dfm[9:0])
      + conv_u2u_10_11(regs_regs_0_1_lpi_3_dfm[19:10])) + conv_u2u_10_12(regs_regs_0_1_lpi_3_dfm[29:20]);
  assign FRAME_acc_6_psp_sva = nl_FRAME_acc_6_psp_sva[11:0];
  assign nl_acc_imod_1_sva = conv_s2s_2_3(conv_s2s_1_2(acc_1_psp_sva[1]) + conv_u2s_1_2(acc_1_psp_sva[0]))
      + conv_s2s_2_3(acc_1_psp_sva[3:2]);
  assign acc_imod_1_sva = nl_acc_imod_1_sva[2:0];
  assign nl_acc_1_psp_sva = (readslicef_5_4_1((conv_u2u_4_5({(readslicef_4_3_1((conv_u2u_3_4({(readslicef_3_2_1((conv_u2u_2_3({(~
      (FRAME_acc_6_psp_sva[3])) , 1'b1}) + conv_u2u_2_3({(FRAME_acc_6_psp_sva[4])
      , (FRAME_acc_6_psp_sva[8])})))) , 1'b1}) + conv_u2u_3_4({(readslicef_3_2_1((conv_u2u_2_3({(~
      (FRAME_acc_6_psp_sva[5])) , 1'b1}) + conv_u2u_2_3({(FRAME_acc_6_psp_sva[6])
      , (~ (FRAME_acc_6_psp_sva[7]))})))) , (FRAME_acc_6_psp_sva[10])})))) , 1'b1})
      + conv_u2u_3_5({(readslicef_3_2_1((conv_u2u_2_3({(~ (FRAME_acc_6_psp_sva[1]))
      , 1'b1}) + conv_u2u_2_3({(FRAME_acc_6_psp_sva[2]) , (~ (FRAME_acc_6_psp_sva[9]))}))))
      , (~ (FRAME_acc_6_psp_sva[11]))})))) + ({3'b101 , (FRAME_acc_6_psp_sva[0])});
  assign acc_1_psp_sva = nl_acc_1_psp_sva[3:0];
  assign and_13_cse = (~(equal_tmp_2 | equal_tmp_1)) & (~(equal_tmp | equal_tmp_3));
  always @(posedge clk) begin
    if ( rst ) begin
      FRAME_p_1_sva <= 3'b0;
      io_read_vout_rsc_d_sdt_1_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg1_lpi_2 <= 6'b0;
      io_read_vout_rsc_d_sdt_sg2_lpi_2 <= 4'b0;
      io_read_vout_rsc_d_sdt_sg3_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg4_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg5_lpi_2 <= 6'b0;
      io_read_vout_rsc_d_sdt_sg6_lpi_2 <= 4'b0;
      io_read_vout_rsc_d_sdt_sg7_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg8_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg9_lpi_2 <= 6'b0;
      io_read_vout_rsc_d_sdt_sg10_lpi_2 <= 4'b0;
      io_read_vout_rsc_d_sdt_sg11_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg12_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg13_lpi_2 <= 6'b0;
      io_read_vout_rsc_d_sdt_sg14_lpi_2 <= 4'b0;
      io_read_vout_rsc_d_sdt_sg15_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg16_lpi_2 <= 10'b0;
      io_read_vout_rsc_d_sdt_sg17_lpi_2 <= 6'b0;
      io_read_vout_rsc_d_sdt_sg18_lpi_2 <= 4'b0;
      io_read_vout_rsc_d_sdt_sg19_lpi_2 <= 10'b0;
      vout_rsc_mgc_out_stdreg_d <= 150'b0;
      SHIFT_i_1_sva_2_sg1 <= 1'b0;
      SHIFT_i_1_sva_3 <= 2'b0;
      regs_regs_0_1_lpi_3 <= 30'b0;
      regs_regs_0_1_lpi_2 <= 30'b0;
      regs_operator_din_1_sva <= 30'b0;
      equal_tmp <= 1'b0;
      equal_tmp_1 <= 1'b0;
      equal_tmp_2 <= 1'b0;
      equal_tmp_3 <= 1'b0;
      regs_regs_0_1_lpi_3_dfm <= 30'b0;
      FRAME_slc_itm <= 1'b0;
      FRAME_p_1_sva_1 <= 3'b0;
      io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm <= 4'b0;
      io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm <= 6'b0;
      io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm <= 4'b0;
      io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm <= 6'b0;
      io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm <= 4'b0;
      io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm <= 6'b0;
      io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm <= 4'b0;
      io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm <= 6'b0;
      io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm <= 10'b0;
      io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm <= 4'b0;
      io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm <= 6'b0;
      io_read_vout_rsc_d_sdt_1_lpi_2_dfm <= 10'b0;
    end
    else begin
      FRAME_p_1_sva <= (MUX_v_3_2_2({FRAME_p_1_sva_1 , FRAME_p_1_sva}, ~((fsm_output[4])
          | (fsm_output[0])))) & (signext_3_1(~ (fsm_output[0])));
      io_read_vout_rsc_d_sdt_1_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_1_lpi_2
          , io_read_vout_rsc_d_sdt_1_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg1_lpi_2 <= MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg1_lpi_2
          , io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg2_lpi_2 <= MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg2_lpi_2
          , io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg3_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg3_lpi_2
          , io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg4_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg4_lpi_2
          , io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg5_lpi_2 <= MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg5_lpi_2
          , io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg6_lpi_2 <= MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg6_lpi_2
          , io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg7_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg7_lpi_2
          , io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg8_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg8_lpi_2
          , io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg9_lpi_2 <= MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg9_lpi_2
          , io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg10_lpi_2 <= MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg10_lpi_2
          , io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg11_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg11_lpi_2
          , io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg12_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg12_lpi_2
          , io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg13_lpi_2 <= MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg13_lpi_2
          , io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg14_lpi_2 <= MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg14_lpi_2
          , io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg15_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg15_lpi_2
          , io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg16_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg16_lpi_2
          , io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg17_lpi_2 <= MUX_v_6_2_2({io_read_vout_rsc_d_sdt_sg17_lpi_2
          , io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg18_lpi_2 <= MUX_v_4_2_2({io_read_vout_rsc_d_sdt_sg18_lpi_2
          , io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm}, fsm_output[4]);
      io_read_vout_rsc_d_sdt_sg19_lpi_2 <= MUX_v_10_2_2({io_read_vout_rsc_d_sdt_sg19_lpi_2
          , io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm}, fsm_output[4]);
      vout_rsc_mgc_out_stdreg_d <= MUX_v_150_2_2({vout_rsc_mgc_out_stdreg_d , ({io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm_mx0 , io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm_mx0
          , io_read_vout_rsc_d_sdt_1_lpi_2_dfm_mx0})}, fsm_output[3]);
      SHIFT_i_1_sva_2_sg1 <= ~ (fsm_output[2]);
      SHIFT_i_1_sva_3 <= (z_out[1:0]) & (signext_2_1(fsm_output[2]));
      regs_regs_0_1_lpi_3 <= MUX1HOT_v_30_4_2({regs_regs_0_1_lpi_2 , regs_operator_din_1_sva
          , regs_regs_0_1_lpi_3 , regs_regs_0_1_lpi_3_dfm}, {(fsm_output[0]) , and_cse
          , (and_34_cse | (~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[0]))))
          , (fsm_output[4])});
      regs_regs_0_1_lpi_2 <= regs_regs_0_1_lpi_3_dfm;
      regs_operator_din_1_sva <= MUX1HOT_v_30_6_2({(vin_rsc_mgc_in_wire_d[29:0])
          , (vin_rsc_mgc_in_wire_d[179:150]) , (vin_rsc_mgc_in_wire_d[329:300]) ,
          (vin_rsc_mgc_in_wire_d[479:450]) , (vin_rsc_mgc_in_wire_d[629:600]) , regs_operator_din_1_sva},
          {(~((FRAME_p_1_sva[2]) | (FRAME_p_1_sva[1]) | (FRAME_p_1_sva[0]) | (fsm_output[2])))
          , ((FRAME_p_1_sva[0]) & nor_7_cse & (~ (fsm_output[2]))) , ((FRAME_p_1_sva[1])
          & nor_8_cse & (~ (fsm_output[2]))) , ((FRAME_p_1_sva[1]) & (FRAME_p_1_sva[0])
          & (~ (FRAME_p_1_sva[2])) & (~ (fsm_output[2]))) , ((FRAME_p_1_sva[2]) &
          nor_9_cse & (~ (fsm_output[2]))) , (fsm_output[2])});
      equal_tmp <= (FRAME_p_1_sva[0]) & nor_7_cse;
      equal_tmp_1 <= (FRAME_p_1_sva[1]) & nor_8_cse;
      equal_tmp_2 <= (FRAME_p_1_sva[1]) & (FRAME_p_1_sva[0]) & (~ (FRAME_p_1_sva[2]));
      equal_tmp_3 <= (FRAME_p_1_sva[2]) & nor_9_cse;
      regs_regs_0_1_lpi_3_dfm <= MUX1HOT_v_30_3_2({regs_regs_0_1_lpi_3_dfm , regs_operator_din_1_sva
          , regs_regs_0_1_lpi_3}, {(~ (fsm_output[2])) , and_cse , and_34_cse});
      FRAME_slc_itm <= readslicef_3_1_2(((z_out[2:0]) + 3'b11));
      FRAME_p_1_sva_1 <= z_out[2:0];
      io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg19_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg18_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg17_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg16_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg15_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg14_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg13_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg12_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg11_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg10_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg9_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg8_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg7_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg6_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg5_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg4_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg3_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg2_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm <= io_read_vout_rsc_d_sdt_sg1_lpi_2_dfm_mx0;
      io_read_vout_rsc_d_sdt_1_lpi_2_dfm <= io_read_vout_rsc_d_sdt_1_lpi_2_dfm_mx0;
    end
  end
  assign mux_47_nl = MUX_v_3_2_2({({SHIFT_i_1_sva_2_sg1 , SHIFT_i_1_sva_3}) , FRAME_p_1_sva},
      fsm_output[3]);
  assign nl_z_out = conv_u2u_3_4(mux_47_nl) + conv_s2u_2_4({(fsm_output[2]) , 1'b1});
  assign z_out = nl_z_out[3:0];

  function [9:0] MUX_v_10_2_2;
    input [19:0] inputs;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[19:10];
      end
      1'b1 : begin
        result = inputs[9:0];
      end
      default : begin
        result = inputs[19:10];
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [3:0] MUX_v_4_2_2;
    input [7:0] inputs;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[7:4];
      end
      1'b1 : begin
        result = inputs[3:0];
      end
      default : begin
        result = inputs[7:4];
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [11:0] inputs;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[11:6];
      end
      1'b1 : begin
        result = inputs[5:0];
      end
      default : begin
        result = inputs[11:6];
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction


  function [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function [5:0] readslicef_7_6_1;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_7_6_1 = tmp[5:0];
  end
  endfunction


  function [3:0] readslicef_5_4_1;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_5_4_1 = tmp[3:0];
  end
  endfunction


  function [2:0] readslicef_4_3_1;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_4_3_1 = tmp[2:0];
  end
  endfunction


  function [5:0] signext_6_2;
    input [1:0] vector;
  begin
    signext_6_2= {{4{vector[1]}}, vector};
  end
  endfunction


  function [1:0] readslicef_3_2_1;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_3_2_1 = tmp[1:0];
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [5:0] inputs;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[5:3];
      end
      1'b1 : begin
        result = inputs[2:0];
      end
      default : begin
        result = inputs[5:3];
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function [149:0] MUX_v_150_2_2;
    input [299:0] inputs;
    input [0:0] sel;
    reg [149:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[299:150];
      end
      1'b1 : begin
        result = inputs[149:0];
      end
      default : begin
        result = inputs[299:150];
      end
    endcase
    MUX_v_150_2_2 = result;
  end
  endfunction


  function [29:0] MUX1HOT_v_30_4_2;
    input [119:0] inputs;
    input [3:0] sel;
    reg [29:0] result;
    integer i;
  begin
    result = inputs[0+:30] & {30{sel[0]}};
    for( i = 1; i < 4; i = i + 1 )
      result = result | (inputs[i*30+:30] & {30{sel[i]}});
    MUX1HOT_v_30_4_2 = result;
  end
  endfunction


  function [29:0] MUX1HOT_v_30_6_2;
    input [179:0] inputs;
    input [5:0] sel;
    reg [29:0] result;
    integer i;
  begin
    result = inputs[0+:30] & {30{sel[0]}};
    for( i = 1; i < 6; i = i + 1 )
      result = result | (inputs[i*30+:30] & {30{sel[i]}});
    MUX1HOT_v_30_6_2 = result;
  end
  endfunction


  function [29:0] MUX1HOT_v_30_3_2;
    input [89:0] inputs;
    input [2:0] sel;
    reg [29:0] result;
    integer i;
  begin
    result = inputs[0+:30] & {30{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*30+:30] & {30{sel[i]}});
    MUX1HOT_v_30_3_2 = result;
  end
  endfunction


  function signed [11:0] conv_u2s_10_12 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_12 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function  [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function  [7:0] conv_u2u_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function signed [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 = {1'b0, vector};
  end
  endfunction


  function signed [11:0] conv_s2s_10_12 ;
    input signed [9:0]  vector ;
  begin
    conv_s2s_10_12 = {{2{vector[9]}}, vector};
  end
  endfunction


  function signed [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 = {1'b0, vector};
  end
  endfunction


  function signed [9:0] conv_s2s_8_10 ;
    input signed [7:0]  vector ;
  begin
    conv_s2s_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function signed [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 = {1'b0, vector};
  end
  endfunction


  function signed [8:0] conv_s2s_7_9 ;
    input signed [6:0]  vector ;
  begin
    conv_s2s_7_9 = {{2{vector[6]}}, vector};
  end
  endfunction


  function signed [6:0] conv_s2s_5_7 ;
    input signed [4:0]  vector ;
  begin
    conv_s2s_5_7 = {{2{vector[4]}}, vector};
  end
  endfunction


  function signed [4:0] conv_s2s_4_5 ;
    input signed [3:0]  vector ;
  begin
    conv_s2s_4_5 = {vector[3], vector};
  end
  endfunction


  function signed [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 = {1'b0, vector};
  end
  endfunction


  function signed [3:0] conv_s2s_3_4 ;
    input signed [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function signed [4:0] conv_s2s_3_5 ;
    input signed [2:0]  vector ;
  begin
    conv_s2s_3_5 = {{2{vector[2]}}, vector};
  end
  endfunction


  function signed [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction


  function  [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function  [11:0] conv_u2u_10_12 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_12 = {{2{1'b0}}, vector};
  end
  endfunction


  function signed [2:0] conv_s2s_2_3 ;
    input signed [1:0]  vector ;
  begin
    conv_s2s_2_3 = {vector[1], vector};
  end
  endfunction


  function signed [1:0] conv_s2s_1_2 ;
    input signed [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function signed [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 = {1'b0, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function  [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [4:0] conv_u2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_5 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [3:0] conv_s2u_2_4 ;
    input signed [1:0]  vector ;
  begin
    conv_s2u_2_4 = {{2{vector[1]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    mean_vga
//  Generated from file(s):
//    2) $PROJECT_HOME/../../../../catapult_proj/vga_blur/blur.c
// ------------------------------------------------------------------


module mean_vga (
  vin_rsc_z, vout_rsc_z, clk, rst
);
  input [749:0] vin_rsc_z;
  output [149:0] vout_rsc_z;
  input clk;
  input rst;


  // Interconnect Declarations
  wire [749:0] vin_rsc_mgc_in_wire_d;
  wire [149:0] vout_rsc_mgc_out_stdreg_d;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire #(.rscid(1),
  .width(750)) vin_rsc_mgc_in_wire (
      .d(vin_rsc_mgc_in_wire_d),
      .z(vin_rsc_z)
    );
  mgc_out_stdreg #(.rscid(2),
  .width(150)) vout_rsc_mgc_out_stdreg (
      .d(vout_rsc_mgc_out_stdreg_d),
      .z(vout_rsc_z)
    );
  mean_vga_core mean_vga_core_inst (
      .clk(clk),
      .rst(rst),
      .vin_rsc_mgc_in_wire_d(vin_rsc_mgc_in_wire_d),
      .vout_rsc_mgc_out_stdreg_d(vout_rsc_mgc_out_stdreg_d)
    );
endmodule



